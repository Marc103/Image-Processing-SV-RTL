package golden_models_pkg;
    import testbench_common_pkg::*;
    import testbench_util_pkg::*;
    import triggerable_queue_pkg::*;
    import camera_simulation_pkg::*;
    import pixel_data_interface_utils_pkg::*;

    `include "util/golden_models/bilinear_xform_model.sv"
    `include "util/golden_models/convolution_model.sv"
    `include "util/golden_models/divisor_model.sv"
    
endpackage