`ifndef _TESTBENCH_UTIL_PKG_SVH
`define _TESTBENCH_UTIL_PKG_SVH

interface clocked_valid_interface (
    input clk,
    input valid
);
endinterface

`endif
